module immediate_generator (