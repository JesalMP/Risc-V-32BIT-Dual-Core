module EX (
    input logic clk,
    input logic rst_n,
    input
    
);
  // EX stage implementation would go here